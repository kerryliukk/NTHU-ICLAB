module pw2num(
    input [8-1:0] pw, 
    output reg [8-1:0] num
);

always @* begin
    case (pw)
        8'd0: num = 8'd1;
        8'd1: num = 8'd2;
        8'd2: num = 8'd4;
        8'd3: num = 8'd8;
        8'd4: num = 8'd16;
        8'd5: num = 8'd32;
        8'd6: num = 8'd64;
        8'd7: num = 8'd128;
        8'd8: num = 8'd29;
        8'd9: num = 8'd58;
        8'd10: num = 8'd116;
        8'd11: num = 8'd232;
        8'd12: num = 8'd205;
        8'd13: num = 8'd135;
        8'd14: num = 8'd19;
        8'd15: num = 8'd38;
        8'd16: num = 8'd76;
        8'd17: num = 8'd152;
        8'd18: num = 8'd45;
        8'd19: num = 8'd90;
        8'd20: num = 8'd180;
        8'd21: num = 8'd117;
        8'd22: num = 8'd234;
        8'd23: num = 8'd201;
        8'd24: num = 8'd143;
        8'd25: num = 8'd3;
        8'd26: num = 8'd6;
        8'd27: num = 8'd12;
        8'd28: num = 8'd24;
        8'd29: num = 8'd48;
        8'd30: num = 8'd96;
        8'd31: num = 8'd192;
        8'd32: num = 8'd157;
        8'd33: num = 8'd39;
        8'd34: num = 8'd78;
        8'd35: num = 8'd156;
        8'd36: num = 8'd37;
        8'd37: num = 8'd74;
        8'd38: num = 8'd148;
        8'd39: num = 8'd53;
        8'd40: num = 8'd106;
        8'd41: num = 8'd212;
        8'd42: num = 8'd181;
        8'd43: num = 8'd119;
        8'd44: num = 8'd238;
        8'd45: num = 8'd193;
        8'd46: num = 8'd159;
        8'd47: num = 8'd35;
        8'd48: num = 8'd70;
        8'd49: num = 8'd140;
        8'd50: num = 8'd5;
        8'd51: num = 8'd10;
        8'd52: num = 8'd20;
        8'd53: num = 8'd40;
        8'd54: num = 8'd80;
        8'd55: num = 8'd160;
        8'd56: num = 8'd93;
        8'd57: num = 8'd186;
        8'd58: num = 8'd105;
        8'd59: num = 8'd210;
        8'd60: num = 8'd185;
        8'd61: num = 8'd111;
        8'd62: num = 8'd222;
        8'd63: num = 8'd161;
        8'd64: num = 8'd95;
        8'd65: num = 8'd190;
        8'd66: num = 8'd97;
        8'd67: num = 8'd194;
        8'd68: num = 8'd153;
        8'd69: num = 8'd47;
        8'd70: num = 8'd94;
        8'd71: num = 8'd188;
        8'd72: num = 8'd101;
        8'd73: num = 8'd202;
        8'd74: num = 8'd137;
        8'd75: num = 8'd15;
        8'd76: num = 8'd30;
        8'd77: num = 8'd60;
        8'd78: num = 8'd120;
        8'd79: num = 8'd240;
        8'd80: num = 8'd253;
        8'd81: num = 8'd231;
        8'd82: num = 8'd211;
        8'd83: num = 8'd187;
        8'd84: num = 8'd107;
        8'd85: num = 8'd214;
        8'd86: num = 8'd177;
        8'd87: num = 8'd127;
        8'd88: num = 8'd254;
        8'd89: num = 8'd225;
        8'd90: num = 8'd223;
        8'd91: num = 8'd163;
        8'd92: num = 8'd91;
        8'd93: num = 8'd182;
        8'd94: num = 8'd113;
        8'd95: num = 8'd226;
        8'd96: num = 8'd217;
        8'd97: num = 8'd175;
        8'd98: num = 8'd67;
        8'd99: num = 8'd134;
        8'd100: num = 8'd17;
        8'd101: num = 8'd34;
        8'd102: num = 8'd68;
        8'd103: num = 8'd136;
        8'd104: num = 8'd13;
        8'd105: num = 8'd26;
        8'd106: num = 8'd52;
        8'd107: num = 8'd104;
        8'd108: num = 8'd208;
        8'd109: num = 8'd189;
        8'd110: num = 8'd103;
        8'd111: num = 8'd206;
        8'd112: num = 8'd129;
        8'd113: num = 8'd31;
        8'd114: num = 8'd62;
        8'd115: num = 8'd124;
        8'd116: num = 8'd248;
        8'd117: num = 8'd237;
        8'd118: num = 8'd199;
        8'd119: num = 8'd147;
        8'd120: num = 8'd59;
        8'd121: num = 8'd118;
        8'd122: num = 8'd236;
        8'd123: num = 8'd197;
        8'd124: num = 8'd151;
        8'd125: num = 8'd51;
        8'd126: num = 8'd102;
        8'd127: num = 8'd204;
        8'd128: num = 8'd133;
        8'd129: num = 8'd23;
        8'd130: num = 8'd46;
        8'd131: num = 8'd92;
        8'd132: num = 8'd184;
        8'd133: num = 8'd109;
        8'd134: num = 8'd218;
        8'd135: num = 8'd169;
        8'd136: num = 8'd79;
        8'd137: num = 8'd158;
        8'd138: num = 8'd33;
        8'd139: num = 8'd66;
        8'd140: num = 8'd132;
        8'd141: num = 8'd21;
        8'd142: num = 8'd42;
        8'd143: num = 8'd84;
        8'd144: num = 8'd168;
        8'd145: num = 8'd77;
        8'd146: num = 8'd154;
        8'd147: num = 8'd41;
        8'd148: num = 8'd82;
        8'd149: num = 8'd164;
        8'd150: num = 8'd85;
        8'd151: num = 8'd170;
        8'd152: num = 8'd73;
        8'd153: num = 8'd146;
        8'd154: num = 8'd57;
        8'd155: num = 8'd114;
        8'd156: num = 8'd228;
        8'd157: num = 8'd213;
        8'd158: num = 8'd183;
        8'd159: num = 8'd115;
        8'd160: num = 8'd230;
        8'd161: num = 8'd209;
        8'd162: num = 8'd191;
        8'd163: num = 8'd99;
        8'd164: num = 8'd198;
        8'd165: num = 8'd145;
        8'd166: num = 8'd63;
        8'd167: num = 8'd126;
        8'd168: num = 8'd252;
        8'd169: num = 8'd229;
        8'd170: num = 8'd215;
        8'd171: num = 8'd179;
        8'd172: num = 8'd123;
        8'd173: num = 8'd246;
        8'd174: num = 8'd241;
        8'd175: num = 8'd255;
        8'd176: num = 8'd227;
        8'd177: num = 8'd219;
        8'd178: num = 8'd171;
        8'd179: num = 8'd75;
        8'd180: num = 8'd150;
        8'd181: num = 8'd49;
        8'd182: num = 8'd98;
        8'd183: num = 8'd196;
        8'd184: num = 8'd149;
        8'd185: num = 8'd55;
        8'd186: num = 8'd110;
        8'd187: num = 8'd220;
        8'd188: num = 8'd165;
        8'd189: num = 8'd87;
        8'd190: num = 8'd174;
        8'd191: num = 8'd65;
        8'd192: num = 8'd130;
        8'd193: num = 8'd25;
        8'd194: num = 8'd50;
        8'd195: num = 8'd100;
        8'd196: num = 8'd200;
        8'd197: num = 8'd141;
        8'd198: num = 8'd7;
        8'd199: num = 8'd14;
        8'd200: num = 8'd28;
        8'd201: num = 8'd56;
        8'd202: num = 8'd112;
        8'd203: num = 8'd224;
        8'd204: num = 8'd221;
        8'd205: num = 8'd167;
        8'd206: num = 8'd83;
        8'd207: num = 8'd166;
        8'd208: num = 8'd81;
        8'd209: num = 8'd162;
        8'd210: num = 8'd89;
        8'd211: num = 8'd178;
        8'd212: num = 8'd121;
        8'd213: num = 8'd242;
        8'd214: num = 8'd249;
        8'd215: num = 8'd239;
        8'd216: num = 8'd195;
        8'd217: num = 8'd155;
        8'd218: num = 8'd43;
        8'd219: num = 8'd86;
        8'd220: num = 8'd172;
        8'd221: num = 8'd69;
        8'd222: num = 8'd138;
        8'd223: num = 8'd9;
        8'd224: num = 8'd18;
        8'd225: num = 8'd36;
        8'd226: num = 8'd72;
        8'd227: num = 8'd144;
        8'd228: num = 8'd61;
        8'd229: num = 8'd122;
        8'd230: num = 8'd244;
        8'd231: num = 8'd245;
        8'd232: num = 8'd247;
        8'd233: num = 8'd243;
        8'd234: num = 8'd251;
        8'd235: num = 8'd235;
        8'd236: num = 8'd203;
        8'd237: num = 8'd139;
        8'd238: num = 8'd11;
        8'd239: num = 8'd22;
        8'd240: num = 8'd44;
        8'd241: num = 8'd88;
        8'd242: num = 8'd176;
        8'd243: num = 8'd125;
        8'd244: num = 8'd250;
        8'd245: num = 8'd233;
        8'd246: num = 8'd207;
        8'd247: num = 8'd131;
        8'd248: num = 8'd27;
        8'd249: num = 8'd54;
        8'd250: num = 8'd108;
        8'd251: num = 8'd216;
        8'd252: num = 8'd173;
        8'd253: num = 8'd71;
        8'd254: num = 8'd142;
        8'd255: num = 8'd1;
        default: num = 8'd0;
    endcase
end

endmodule